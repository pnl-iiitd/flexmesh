
wire kernel_monitor_reset;
wire kernel_monitor_clock;
wire kernel_monitor_report;
assign kernel_monitor_reset = ~ap_rst_n;
assign kernel_monitor_clock = ap_clk;
assign kernel_monitor_report = 1'b0;
wire [6:0] axis_block_sigs;
wire [6:0] inst_idle_sigs;
wire [0:0] inst_block_sigs;
wire kernel_block;

assign axis_block_sigs[0] = ~out_s_TDATA_blk_n;
assign axis_block_sigs[1] = ~grp_read_stream_fu_1501.in_s_TDATA_blk_n;
assign axis_block_sigs[2] = ~grp_read_stream_fu_1501.grp_read_stream_Pipeline_IV_stream_read_fu_168.in_s_TDATA_blk_n;
assign axis_block_sigs[3] = ~grp_read_stream_fu_1501.grp_read_stream_Pipeline_PT_stream_read_fu_189.in_s_TDATA_blk_n;
assign axis_block_sigs[4] = ~grp_read_stream_fu_1501.grp_read_stream_Pipeline_AAD_stream_read_fu_204.in_s_TDATA_blk_n;
assign axis_block_sigs[5] = ~grp_read_stream_fu_1501.grp_read_stream_Pipeline_Key_stream_read_fu_221.in_s_TDATA_blk_n;
assign axis_block_sigs[6] = ~grp_GCM_AE_HW_1x1_Pipeline_cipher_text_array_to_stream_fu_2323.out_s_TDATA_blk_n;

assign inst_block_sigs[0] = 1'b0;

assign inst_idle_sigs[0] = 1'b0;
assign inst_idle_sigs[1] = grp_read_stream_fu_1501.ap_idle;
assign inst_idle_sigs[2] = grp_read_stream_fu_1501.grp_read_stream_Pipeline_IV_stream_read_fu_168.ap_idle;
assign inst_idle_sigs[3] = grp_read_stream_fu_1501.grp_read_stream_Pipeline_PT_stream_read_fu_189.ap_idle;
assign inst_idle_sigs[4] = grp_read_stream_fu_1501.grp_read_stream_Pipeline_AAD_stream_read_fu_204.ap_idle;
assign inst_idle_sigs[5] = grp_read_stream_fu_1501.grp_read_stream_Pipeline_Key_stream_read_fu_221.ap_idle;
assign inst_idle_sigs[6] = grp_GCM_AE_HW_1x1_Pipeline_cipher_text_array_to_stream_fu_2323.ap_idle;

GCM_AE_HW_1x1_hls_deadlock_idx0_monitor GCM_AE_HW_1x1_hls_deadlock_idx0_monitor_U (
    .clock(kernel_monitor_clock),
    .reset(kernel_monitor_reset),
    .axis_block_sigs(axis_block_sigs),
    .inst_idle_sigs(inst_idle_sigs),
    .inst_block_sigs(inst_block_sigs),
    .block(kernel_block)
);


always @ (kernel_block or kernel_monitor_reset) begin
    if (kernel_block == 1'b1 && kernel_monitor_reset == 1'b0) begin
        find_kernel_block = 1'b1;
    end
    else begin
        find_kernel_block = 1'b0;
    end
end
